-- -------------------------------------------------------------
-- 
-- Module: MATRIX
-- 
-- -------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.work_pack.all;

entity MATRIX_CTRL is
  generic (
    N  : integer := 50;
    BW : integer := 8
  );
  port( clk						:   in    std_logic;
        reset					:   in    std_logic;
        clk_enable				:   in    std_logic;
        PHASE_in				:   in    std_logic_vector(7 downto 0);  -- int8
        ce_out					:   out   std_logic;
        CONTROL_COEFF			:   out   std_logic_vector(7 downto 0);  -- int8
	    COUNTER_FLAG			:   out   std_logic;
	     
	    wvalid                : in std_logic;
	    wcoladdr              : in unsigned(11 downto 0);
	    wdata                 : in std_logic_vector(N * BW - 1 downto 0)
  );
end MATRIX_CTRL;


architecture rtl of MATRIX_CTRL is

  constant Stages : integer := 3;
  
  signal valid, first : std_logic_vector(Stages - 1 downto 0); 

  -- signals
  signal PHASE_in_signed, inp_ff1, inp_ff2, inp_ff3	: signed(7 downto 0);  -- int8
  signal PHASE_in_unsigned					: unsigned(7 downto 0);  -- int8
  
  signal accum : vector_of_signed8(0 to N - 1);
  
  signal CONTROL_COEFF_array				: vector_of_signed8(0 to N-1);
  signal CONTROL_COEFF_array_final			: vector_of_signed8(0 to N-1);
  signal CONTROL_COEFF_array_final_loop	: vector_of_signed8(0 to N-1);
  
  signal CTRL_unsigned								: unsigned(11 downto 0);  -- int8
  
  signal Multiport_Switch_out				: signed(7 downto 0);  -- int8
  
  signal switch_compare						: std_logic;  -- boolean
  signal ce										: std_logic;  -- boolean
  
  signal counter_up							: unsigned(11 downto 0) := X"fff";
  
  signal koeff_ff1, koeff_ff2, koeff_ff3 : std_logic_vector((N) * BW - 1 downto 0); 
  
  type matrix is array(natural range <>) of std_logic_vector(N * BW - 1 downto 0);

  signal Jij : matrix(0 to N-1);
  constant Jinit : memory := (											
    ('0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('1','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('1','1','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','1','0','0','0','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','1','0','0','0','1','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','1','0','0','0','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','1','0','0','1','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','1','0','0','0','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','1','0','0','0','1','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','1','0','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','1','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
    ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')	);
    
begin


	PHASE_in_signed <= to_signed(1, PHASE_in_signed'length)		 when to_integer(unsigned(PHASE_in(7 downto 0))) >= to_unsigned(16#90#, 8) else
							 to_signed(-1, PHASE_in_signed'length)    when to_integer(unsigned(PHASE_in(7 downto 0))) <= to_unsigned(16#8E#, 8) else
							 to_signed(0, PHASE_in_signed'length);


  ce <= '1';
  
    
  CONTROL_COEFF_array <= accum;         
  
  process (clk, reset)
  variable product : signed(15 downto 0);
  variable col, rev_row : integer;
  variable one_row : std_logic_vector(N * BW - 1 downto 0);
  variable valid_now, first_now : std_logic;
  begin
    if (reset = '1') then
      accum <= (others => (others => '0'));
      valid <= (others => '0');
      first <= (others => '0');
      for row in 0 to N - 1 loop
        for col in 0 to N - 1 loop 
          if Jinit(row, N - 1 - col) = '1' then 
            one_row((col + 1) * BW - 1 downto col * BW) := X"01";
          else 
            one_row((col + 1) * BW - 1 downto col * BW) := X"00";
          end if; 
        end loop; 
        Jij(row) <= one_row;
      end loop; 
    elsif clk'event and clk = '1' then      
      col := to_integer(counter_up);
      if col < N then 
        valid_now := '1';
      else
        valid_now := '0';
      end if;
      
      if col = 0 then
        first_now := '1';
      else
        first_now := '0';
      end if;
      
      inp_ff3 <= inp_ff2;
      inp_ff2 <= inp_ff1;
      inp_ff1 <= PHASE_in_signed;
      
            -- the matrix is turned over a bit, because original code turned over the input vector
      if valid_now = '1' then 
        koeff_ff1 <= Jij(N - 1 - col);
      end if; 
      koeff_ff3 <= koeff_ff2;
      koeff_ff2 <= koeff_ff1;
      
      valid <= valid(Stages - 2 downto 0) & valid_now;
      first <= first(Stages - 2 downto 0) & first_now;
      
      if valid(2) = '1' then
          for row in 0 to N - 1 loop
            rev_row := N - 1 - row;
            product := inp_ff3 * signed(koeff_ff3((rev_row + 1) * BW - 1 downto rev_row * BW));
            if first(2) = '1' then
              accum(row) <= product(7 downto 0);
            else
              accum(row) <= accum(row) + product(7 downto 0);
            end if;
          end loop;
        end if;
    end if;
  end process;
        

  Counter_process : process(clk,reset)
  begin
	if rising_edge(clk) then
		if reset = '1' then
			counter_up <= to_unsigned(16#000#, 12);
		elsif ce = '1' then
			if counter_up < to_unsigned(N + 7, 12) then
				counter_up <= counter_up + 1;
			else 
			counter_up <= to_unsigned(16#00#, 12);
			end if;
		end if;
	end if;
  end process;

  
  Delays2_process : PROCESS (clk, reset)
  BEGIN
    IF reset = '1' THEN
      CONTROL_COEFF_array_final_loop <= (others => to_signed(16#00#, 8));
    ELSIF clk'EVENT AND clk = '1'  THEN
        for i in 0 to N-1 loop 
          CONTROL_COEFF_array_final_loop(i) <= CONTROL_COEFF_array_final(i);
        end loop;
    END IF;
  END PROCESS Delays2_process;  
  
  COUNTER_FLAG <= '1' when counter_up = to_unsigned(16#2B#, 12) else '0';
  
  holdongen: for k in 0 to N-1 generate
  
    CONTROL_COEFF_array_final(k) <= CONTROL_COEFF_array(k) when counter_up = to_unsigned(N + 3, 12) else CONTROL_COEFF_array_final_loop(k);
	
  end generate;
  
  CTRL_unsigned <= counter_up;
  
  Multiport_Switch_out <=
                                CONTROL_COEFF_array_final(N-1 - (TO_INTEGER(CTRL_unsigned) - 16#35#)) when CTRL_unsigned >= to_unsigned(16#35#, 8) and CTRL_unsigned <= to_unsigned(16#39#, 8) else
								CONTROL_COEFF_array_final(44 - (TO_INTEGER(CTRL_unsigned))) when CTRL_unsigned >= to_unsigned(16#0#, 8) and CTRL_unsigned <= to_unsigned(16#2C#, 8) else
								(others => '0');

  CONTROL_COEFF  <= std_logic_vector(Multiport_Switch_out);

  ce_out <= clk_enable;

end rtl;
